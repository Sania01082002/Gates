module or_gate(y,a,b);
input a,b;
output y;
or(y,a,b);
endmodule
